module week0303fi_tb;

reg [3:0] A;
reg [3:0] B;
wire Eq;
wire Gt;
wire Lt;

week0303fi
 U0 (
  .A(A),
  .B(B),
  .Eq(Eq),
  .Gt(Gt),
  .Lt(Lt));

  initial
  begin
    A = 4'b0000;
    #800 A = 4'b0001;
    #800 A = 4'b0010;
    #800 A = 4'b0011;
    #800 A = 4'b0100;
    #800 A = 4'b0101;
    #800 A = 4'b0110;
    #800 A = 4'b0111;
    #800 A = 4'b1000;
    #800 A = 4'b1001;
    #800 A = 4'b1010;
    #800 A = 4'b1011;
    #800 A = 4'b1100;
  end

  initial
  begin
    B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
    #50 B = 4'b1000;
    #50 B = 4'b1001;
    #50 B = 4'b1010;
    #50 B = 4'b1011;
    #50 B = 4'b1100;
    #50 B = 4'b1101;
    #50 B = 4'b1110;
    #50 B = 4'b1111;
    #50 B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
    #50 B = 4'b1000;
    #50 B = 4'b1001;
    #50 B = 4'b1010;
    #50 B = 4'b1011;
    #50 B = 4'b1100;
    #50 B = 4'b1101;
    #50 B = 4'b1110;
    #50 B = 4'b1111;
    #50 B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
    #50 B = 4'b1000;
    #50 B = 4'b1001;
    #50 B = 4'b1010;
    #50 B = 4'b1011;
    #50 B = 4'b1100;
    #50 B = 4'b1101;
    #50 B = 4'b1110;
    #50 B = 4'b1111;
    #50 B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
    #50 B = 4'b1000;
    #50 B = 4'b1001;
    #50 B = 4'b1010;
    #50 B = 4'b1011;
    #50 B = 4'b1100;
    #50 B = 4'b1101;
    #50 B = 4'b1110;
    #50 B = 4'b1111;
    #50 B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
    #50 B = 4'b1000;
    #50 B = 4'b1001;
    #50 B = 4'b1010;
    #50 B = 4'b1011;
    #50 B = 4'b1100;
    #50 B = 4'b1101;
    #50 B = 4'b1110;
    #50 B = 4'b1111;
    #50 B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
    #50 B = 4'b1000;
    #50 B = 4'b1001;
    #50 B = 4'b1010;
    #50 B = 4'b1011;
    #50 B = 4'b1100;
    #50 B = 4'b1101;
    #50 B = 4'b1110;
    #50 B = 4'b1111;
    #50 B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
    #50 B = 4'b1000;
    #50 B = 4'b1001;
    #50 B = 4'b1010;
    #50 B = 4'b1011;
    #50 B = 4'b1100;
    #50 B = 4'b1101;
    #50 B = 4'b1110;
    #50 B = 4'b1111;
    #50 B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
    #50 B = 4'b1000;
    #50 B = 4'b1001;
    #50 B = 4'b1010;
    #50 B = 4'b1011;
    #50 B = 4'b1100;
    #50 B = 4'b1101;
    #50 B = 4'b1110;
    #50 B = 4'b1111;
    #50 B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
    #50 B = 4'b1000;
    #50 B = 4'b1001;
    #50 B = 4'b1010;
    #50 B = 4'b1011;
    #50 B = 4'b1100;
    #50 B = 4'b1101;
    #50 B = 4'b1110;
    #50 B = 4'b1111;
    #50 B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
    #50 B = 4'b1000;
    #50 B = 4'b1001;
    #50 B = 4'b1010;
    #50 B = 4'b1011;
    #50 B = 4'b1100;
    #50 B = 4'b1101;
    #50 B = 4'b1110;
    #50 B = 4'b1111;
    #50 B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
    #50 B = 4'b1000;
    #50 B = 4'b1001;
    #50 B = 4'b1010;
    #50 B = 4'b1011;
    #50 B = 4'b1100;
    #50 B = 4'b1101;
    #50 B = 4'b1110;
    #50 B = 4'b1111;
    #50 B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
    #50 B = 4'b1000;
    #50 B = 4'b1001;
    #50 B = 4'b1010;
    #50 B = 4'b1011;
    #50 B = 4'b1100;
    #50 B = 4'b1101;
    #50 B = 4'b1110;
    #50 B = 4'b1111;
    #50 B = 4'b0000;
    #50 B = 4'b0001;
    #50 B = 4'b0010;
    #50 B = 4'b0011;
    #50 B = 4'b0100;
    #50 B = 4'b0101;
    #50 B = 4'b0110;
    #50 B = 4'b0111;
  end

endmodule
