module week02s02_tb;

reg [1:0] A;
reg [1:0] B;
wire Eq;
wire Gt;
wire Lt;

week02s02
 U0 (
  .A(A),
  .B(B),
  .Eq(Eq),
  .Gt(Gt),
  .Lt(Lt));

  initial
  begin
    A = 2'b00;
    #200 A = 2'b01;
    #200 A = 2'b10;
    #200 A = 2'b11;
    #200 A = 2'b00;
    #200 A = 2'b01;
    #200 A = 2'b10;
    #200 A = 2'b11;
    #200 A = 2'b00;
    #200 A = 2'b01;
    #200 A = 2'b10;
    #200 A = 2'b11;
    #200 A = 2'b00;
    #200 A = 2'b01;
    #200 A = 2'b10;
    #200 A = 2'b11;
    #200 A = 2'b00;
    #200 A = 2'b01;
    #200 A = 2'b10;
    #200 A = 2'b11;
    #200 A = 2'b00;
    #200 A = 2'b01;
    #200 A = 2'b10;
    #200 A = 2'b11;
    #200 A = 2'b00;
    #200 A = 2'b01;
    #200 A = 2'b10;
    #200 A = 2'b11;
    #200 A = 2'b00;
    #200 A = 2'b01;
    #200 A = 2'b10;
    #200 A = 2'b11;
    #200 A = 2'b00;
    #200 A = 2'b01;
    #200 A = 2'b10;
    #200 A = 2'b11;
    #200 A = 2'b00;
    #200 A = 2'b01;
    #200 A = 2'b10;
    #200 A = 2'b11;
    #200 A = 2'b00;
    #200 A = 2'b01;
    #200 A = 2'b10;
    #200 A = 2'b11;
    #200 A = 2'b00;
    #200 A = 2'b01;
    #200 A = 2'b10;
    #200 A = 2'b11;
    #200 A = 2'b00;
    #200 A = 2'b01;
  end

  initial
  begin
    B = 2'b00;
    #400 B = 2'b01;
    #400 B = 2'b10;
    #400 B = 2'b11;
    #400 B = 2'b00;
    #400 B = 2'b01;
    #400 B = 2'b10;
    #400 B = 2'b11;
    #400 B = 2'b00;
    #400 B = 2'b01;
    #400 B = 2'b10;
    #400 B = 2'b11;
    #400 B = 2'b00;
    #400 B = 2'b01;
    #400 B = 2'b10;
    #400 B = 2'b11;
    #400 B = 2'b00;
    #400 B = 2'b01;
    #400 B = 2'b10;
    #400 B = 2'b11;
    #400 B = 2'b00;
    #400 B = 2'b01;
    #400 B = 2'b10;
    #400 B = 2'b11;
    #400 B = 2'b00;
  end

endmodule
