module week030201_tb;

reg [9:0] A;
reg [9:0] B;
wire CHK2;
wire [4:0] Sum;

week030201
 U0 (
  .A(A),
  .B(B),
  .CHK2(CHK2),
  .Sum(Sum));

  initial
  begin
    A = 10'b1000000000;
    #2000 A = 10'b0000000000;
    #100 A = 10'b0001000000;
  end

  initial
  begin
    B = 10'b1000000000;
    #100 B = 10'b0100000000;
    #100 B = 10'b0010000000;
    #100 B = 10'b0001000000;
    #100 B = 10'b0000100000;
    #100 B = 10'b0000010000;
    #100 B = 10'b0000001000;
    #100 B = 10'b0000000100;
    #100 B = 10'b0000000010;
    #100 B = 10'b0000000001;
    #100 B = 10'b0000000000;
    #1100 B = 10'b1000000000;
    #100 B = 10'b0000000000;
    #100 B = 10'b0100000000;
    #100 B = 10'b0000000000;
    #100 B = 10'b0010000000;
    #100 B = 10'b0000000000;
    #100 B = 10'b0000001000;
    #100 B = 10'b0000000000;
    #200 B = 10'b0000000010;
    #100 B = 10'b0000000000;
  end

endmodule
